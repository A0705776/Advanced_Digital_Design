module ButtonTest(in,out);
	input in;
	output[6:0] out;
	
	CheckButton(in,out);
	
endmodule
